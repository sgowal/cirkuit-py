innerBorder = 125,253,126,265,137,271,149,271,161,272,174,284,176,304,174,320,174,334,174,349,173,359,161,374,147,374,134,374,125,375,124,385,132,386,147,388,163,390,171,412,170,422,170,443,167,458,167,471,153,483,139,488,120,489,118,500,203,499,207,407,215,394,229,390,243,389,258,385,257,350,257,321,261,315,269,312,269,299,269,284,267,260,267,248,254,233,250,165,246,144,249,126,245,109,131,106
tolerance = 10
name = Challenge
maximumSpeed = 7
startingLine = 67,142,137,142
outerBorder = 97,44,82,63,79,77,79,102,77,287,78,304,86,313,101,314,132,317,135,327,131,336,102,336,84,337,77,345,77,358,77,378,77,394,77,407,85,419,98,420,120,421,130,429,130,440,121,445,107,445,94,445,82,444,73,452,73,467,73,483,73,500,73,515,74,536,92,552,119,554,173,553,214,553,240,554,255,540,257,518,257,503,257,487,257,463,257,449,272,442,293,440,312,438,321,429,321,407,319,381,318,346,317,322,308,315,307,305,307,296,307,283,305,252,312,243,318,236,316,173,314,147,314,131,314,115,314,94,304,71,289,55,272,49,249,44,112,40
