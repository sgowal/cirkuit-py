innerBorder = 506,171,526,205,527,243,513,250,490,248,464,238,432,226,403,222,385,239,373,268,371,294,404,297,445,305,458,331,436,348,391,347,359,351,352,386,362,470,367,512,351,496,340,467,333,445,324,409,306,381,281,364,259,360,251,377,246,402,238,425,224,441,206,445,170,436,149,425,127,396,115,359,124,321,139,302,159,286,177,277,206,265,224,250,229,232,230,214,219,200,206,190,181,180,154,174,122,167,112,154,111,113,120,103,143,91,187,78,217,70,247,68,297,68,337,74,366,81,392,89,417,100,448,117,473,131,487,142
tolerance = 10
name = Complex
maximumSpeed = 8
startingLine = 136,137,30,137
outerBorder = 530,70,560,100,580,149,585,194,583,238,570,272,538,290,477,275,437,263,474,279,501,328,487,390,434,393,396,397,401,442,409,487,407,519,396,543,373,551,343,542,320,520,310,504,296,481,288,441,279,408,272,434,254,490,213,500,183,496,132,481,108,466,86,445,71,423,54,377,59,336,79,304,97,290,124,267,159,237,169,228,155,224,112,217,74,195,50,168,49,112,63,69,96,39,149,24,218,12,255,11,325,11,382,15,438,27,473,37
